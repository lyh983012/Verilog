`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:56:59 06/01/2014 
// Design Name: 
// Module Name:    intel8056 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module intel8056(
    output SA0,SA1,SA2,SA3,SA4,SA5,SA6,SA7,SA8,SA9,
    output IOR,
    output IOW,
    output [7:0] SD,
    inout GND,
    input AEN
    );


endmodule
