`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:11:25 06/01/2014 
// Design Name: 
// Module Name:    my8056 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module my8056(
    output SA0,
    output SA1,
    output SA2,
    output SA3,
    output SA4,
    output SA5,
    output SA6,
    output SA7,
    output SA8,
    output SA9,
    output IOR,
    output IOW,
    output AEN,
    inout GND,
    output [7:0] SD
    );


endmodule
